library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity processador is
    Port (
        
    );
end processador;

architecture Behavioral of processador is

begin



end Behavioral;
